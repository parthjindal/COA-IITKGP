`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:11:34 11/07/2021 
// Design Name: 
// Module Name:    PC 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module PC(
    input [31:0] inp,
	 input clk,
	 input rst,
	 output reg [31:0] out
    );
	 
	 always @(negedge clk or posedge rst) begin
	    if (rst)
		     out <= 10'b0;
		 else out <= inp;
	 end

endmodule
