`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:03:34 11/07/2021 
// Design Name: 
// Module Name:    UpdatePC 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module UpdatePC(
    input [31:0] in,
	 input lblSel,
	 input jumpSel,
	 input branch,
	 input [25:0] label1,
	 input [31:0] label2,
	 output [31:0] 
    );


endmodule
