`timescale 10ns/1ps

module LFSR;
endmodule
