`timescale 1ns/1ps

module booth_multiplier();
  // skeleton
endmodule
