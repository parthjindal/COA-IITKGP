`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Assignment: 05
// Engineeer: Parth Jindal, Pranav Rajput Group 024
// Module Name: MUX 
// Description: 2-1 Multiplexer
//////////////////////////////////////////////////////////////////////////////////
module MUX(
    output Out,
    input d0,
    input d1,
    input sel
    );
	assign Out = (sel) ? d1 : d0;
endmodule
