'timescale 10ns/1ps

module testBench;
endmodule
